* NGSPICE file created from Inverter.ext - technology: sky130B

.subckt sky130_fd_pr__nfet_g5v0d10v5_6XHARQ a_n108_n75# a_n50_n163# a_n242_n297# a_50_n75#
X0 a_50_n75# a_n50_n163# a_n108_n75# a_n242_n297# sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7EBZY6 a_50_n150# a_n50_n247# a_n108_n150# w_n308_n447#
X0 a_50_n150# a_n50_n247# a_n108_n150# w_n308_n447# sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
.ends

.subckt Inverter Vin VDD VSS Vout
XXM1 VSS Vin VSS Vout sky130_fd_pr__nfet_g5v0d10v5_6XHARQ
XXM2 Vout Vin VDD VDD sky130_fd_pr__pfet_g5v0d10v5_7EBZY6
.ends

